
module encoder(
  in,
  out
  );
 
  input wire [7:0] in; 
  output reg [2:0] out;
        
  always @ (*) begin
    casex (in)
      8'b???????1 : out = 0;
      8'b??????1? : out = 1; 
      8'b?????1?? : out = 2; 
      8'b????1??? : out = 3; 
      8'b???1???? : out = 4;
      8'b??1????? : out = 5; 
      8'b?1?????? : out = 6; 
      8'b1??????? : out = 7;
   endcase
  end

endmodule
