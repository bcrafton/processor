`ifndef _defines_vh_
`define _defines_vh_

`define DATA_WIDTH 16

`endif
