
module encoder3x8(
  in,
  out
  );
 
  input wire [7:0] in; 
  output reg [2:0] out;
        
  always @ (*) begin
    casex (in)
      8'b???????1 : out = 0;
      8'b??????1? : out = 1; 
      8'b?????1?? : out = 2; 
      8'b????1??? : out = 3; 
      8'b???1???? : out = 4;
      8'b??1????? : out = 5; 
      8'b?1?????? : out = 6; 
      8'b1??????? : out = 7;
    endcase
  end

endmodule


module encoder5x32(
  in,
  out
  );
 
  input wire [31:0] in; 
  output reg [4:0] out;
        
  always @ (*) begin
    casex (in)
      32'b???????????????????????????????1 : out = 0;
      32'b??????????????????????????????1? : out = 1;
      32'b?????????????????????????????1?? : out = 2;
      32'b????????????????????????????1??? : out = 3;

      32'b???????????????????????????1???? : out = 4;
      32'b??????????????????????????1????? : out = 5;
      32'b?????????????????????????1?????? : out = 6;
      32'b????????????????????????1??????? : out = 7;

      32'b???????????????????????1???????? : out = 8;
      32'b??????????????????????1????????? : out = 9;
      32'b?????????????????????1?????????? : out = 10;
      32'b????????????????????1??????????? : out = 11;

      32'b???????????????????1???????????? : out = 12;
      32'b??????????????????1????????????? : out = 13;
      32'b?????????????????1?????????????? : out = 14;
      32'b????????????????1??????????????? : out = 15;

      32'b???????????????1???????????????? : out = 16;
      32'b??????????????1????????????????? : out = 17;
      32'b?????????????1?????????????????? : out = 18;
      32'b????????????1??????????????????? : out = 19;

      32'b???????????1???????????????????? : out = 20;
      32'b??????????1????????????????????? : out = 21;
      32'b?????????1?????????????????????? : out = 22;
      32'b????????1??????????????????????? : out = 23;

      32'b???????1???????????????????????? : out = 24;
      32'b??????1????????????????????????? : out = 25;
      32'b?????1?????????????????????????? : out = 26;
      32'b????1??????????????????????????? : out = 27;

      32'b???1???????????????????????????? : out = 28;
      32'b??1????????????????????????????? : out = 29;
      32'b?1?????????????????????????????? : out = 30;
      32'b1??????????????????????????????? : out = 31;
    endcase
  end

endmodule
